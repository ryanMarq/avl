../../template/rtl/example_hdl.sv