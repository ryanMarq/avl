module example_hdl();

    logic        clk;
    logic        rst_n;
    logic [31:0] data;

endmodule : example_hdl
